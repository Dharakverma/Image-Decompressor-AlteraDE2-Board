library verilog;
use verilog.vl_types.all;
entity M2_Multiplier is
    port(
        op1             : in     integer;
        op2             : in     integer;
        \out\           : out    integer
    );
end M2_Multiplier;
